// -----------------------------------------------------------------------------
// Copyright (c) 2014-2019 All rights reserved
// -----------------------------------------------------------------------------
// Author : Javen   penguinleo@163.com
// File   : ModelSelModule.v
// Create : 2020-08-11 11:48:15
// Revise : 2020-08-11 11:48:15
// Editor : sublime text3, tab size (4)
// Comment: This module is a logic definition moudle for the UART module work mode select.
//  		different mode value set would make the uart module in normal mode, auto-echo, local loopback
// 			remote looback.
//          Up module:
//              
//          Sub module:
//             
// Input Signal List:
//      1   |   CLK                 :   clock signal
//      2   |   RST                 :   reset signal
//      3   | 
// Output Signal List:      
//      1   |                                                                                             |  
// Note:  
// -----------------------------------------------------------------------------   